`ifndef __l_class_OC_foo_VH__
`define __l_class_OC_foo_VH__

`define l_class_OC_foo_RULE_COUNT (0)

//METAWRITE; indication$heard; :stop_main_program;
//METAGUARD; indication$heard__RDY; 1;
`endif

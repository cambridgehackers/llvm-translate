`ifndef __l_class_OC_Echo_VH__
`define __l_class_OC_Echo_VH__

`define l_class_OC_Echo_RULE_COUNT (0)

//METAINVOKE; request$say; :indication$heard;
//METAGUARD; request$say; indication$heard__RDY;
//METAEXTERNAL; indication; l_class_OC_EchoIndication;
`endif

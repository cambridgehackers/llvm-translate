module top(input CLK, input nRST);
  always @( posedge CLK) begin
    if (!nRST) then begin
    end
    else begin
//processing printf

    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


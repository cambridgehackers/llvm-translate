module l_class_OC_Echo (
    input CLK,
    input nRST);

  ;
  ;
   reg[31:0] pipetemp;
  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


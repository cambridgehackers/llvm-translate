`ifndef __l_class_OC_EchoRequestOutput_VH__
`define __l_class_OC_EchoRequestOutput_VH__

`define l_class_OC_EchoRequestOutput_RULE_COUNT (0)

//METAEXTERNAL; pipe; l_class_OC_PipeIn_OC_0;
`endif

module top(input CLK, input nRST);
  always @( posedge CLK) begin
    if (!nRST) then begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


interface L_class_OC_Echo_KD__KD_respond;
endinterface
import "BVI" l_class_OC_Echo_KD__KD_respond =
module mkL_class_OC_Echo_KD__KD_respond(L_class_OC_Echo_KD__KD_respond);
    default_reset rst(nRST);
    default_clock clk(CLK);
    schedule () CF ();
endmodule

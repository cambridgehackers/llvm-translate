`ifndef __l_class_OC_EchoRequestInput_VH__
`define __l_class_OC_EchoRequestInput_VH__

`define l_class_OC_EchoRequestInput_RULE_COUNT (0)

//METAEXTERNAL; request; l_class_OC_EchoRequest;
//METAREAD; pipe_enq; :;pipe_enq_v$tag:pipe_enq_v$tag == 1;pipe_enq_v$data$say$meth:;pipe_enq_v$tag:pipe_enq_v$tag == 1;pipe_enq_v$data$say$v:;pipe_enq_v$tag;
//METAINVOKE; pipe_enq; :pipe_enq_v$tag == 1;request$say;
//METAGUARD; pipe_enq__RDY; request$say__RDY;
`endif

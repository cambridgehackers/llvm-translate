`ifndef __l_class_OC_Echo_VH__
`define __l_class_OC_Echo_VH__

`define l_class_OC_Echo_RULE_COUNT (0)

//METAEXTERNAL; indication; l_class_OC_EchoIndication;
//METAINVOKE; request$say; :indication$heard;
//METAGUARD; request$say__RDY; indication$heard__RDY;
`endif

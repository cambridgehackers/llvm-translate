module l_class_OC_EchoRequest (
    input CLK,
    input nRST);
    always @( posedge CLK) begin
      if (!nRST) begin
      end // nRST
    end // always @ (posedge CLK)
endmodule 


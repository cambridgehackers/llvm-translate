module l_class_OC_Rule (
    input CLK,
    input nRST);

   reg[31:0]  (**_vptr_EC_Rule) ( VERILOG_int, ...);
  ;
  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


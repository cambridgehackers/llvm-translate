module l_class_OC_Echo_KD__KD_respond (
    input CLK,
    input nRST);

  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


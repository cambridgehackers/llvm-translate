module l_class_OC_Fifo (
    input CLK,
    input nRST);
  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


module l_class_OC_Module (
    input CLK,
    input nRST);

  ;
  ;
  VERILOGunsigned VERILOG_long long size;
  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 


`ifndef __l_class_OC_EchoIndicationOutput_VH__
`define __l_class_OC_EchoIndicationOutput_VH__

`define l_class_OC_EchoIndicationOutput_RULE_COUNT (0)

//METAWRITE; indication$heard; :ind$data$heard$meth;:ind$data$heard$v;
//METAINVOKE; indication$heard; :pipe$enq;
//METAGUARD; indication$heard; pipe$enq__RDY;
//METAEXTERNAL; pipe; l_class_OC_PipeIn_OC_0;
`endif

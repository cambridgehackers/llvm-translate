
//METARULES; A; B; C
//METAGUARD; A__RDY; ACond
//METAGUARD; B__RDY; BCond
//METAGUARD; C__RDY; CCond

//METAWRITE; A; 1; 2; 3
//METAREAD; A; 4; 5; 6
//METAWRITE; B; 6
//METAREAD; B; 4; 7
//METAWRITE; C; 7; 8; 5
//METAREAD; C; 4

`ifndef __l_class_OC_EchoRequestOutput_VH__
`define __l_class_OC_EchoRequestOutput_VH__

`define l_class_OC_EchoRequestOutput_RULE_COUNT (0)

//METAEXTERNAL; pipe; l_class_OC_PipeIn;
//METAGUARD; say__RDY; pipe$enq__RDY;
//METAWRITE; say; :;ind$data$say$meth:;ind$data$say$v;
//METAINVOKE; say; :;pipe$enq;
`endif

interface L_class_OC_EchoRequestOutput;
endinterface
import "BVI" l_class_OC_EchoRequestOutput =
module mkL_class_OC_EchoRequestOutput(L_class_OC_EchoRequestOutput);
    default_reset rst(nRST);
    default_clock clk(CLK);
    schedule () CF ();
endmodule

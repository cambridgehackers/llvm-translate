interface L_class_OC_EchoIndicationOutput;
endinterface
import "BVI" l_class_OC_EchoIndicationOutput =
module mkL_class_OC_EchoIndicationOutput(L_class_OC_EchoIndicationOutput);
    default_reset rst(nRST);
    default_clock clk(CLK);
    schedule () CF ();
endmodule

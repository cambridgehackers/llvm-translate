`ifndef __l_class_OC_EchoRequestOutput_VH__
`define __l_class_OC_EchoRequestOutput_VH__

`define l_class_OC_EchoRequestOutput_RULE_COUNT (0)

//METAEXTERNAL; pipe; l_class_OC_PipeIn;
//METAGUARD; request$say__RDY; pipe$enq__RDY;
//METAWRITE; request$say; :ind$data$say$meth;:ind$data$say$v;
//METAINVOKE; request$say; :pipe$enq;
`endif


//METARULES; A; B; C; E; F
//METAGUARD; A__RDY; ACond
//METAGUARD; B__RDY; BCond
//METAGUARD; C__RDY; CCond
//METAGUARD; D__RDY; DCond
//METAGUARD; E__RDY; ECond
//METAGUARD; F__RDY; FCond

//METAWRITE; B; 6
//METAREAD; B; 4; 7; 9
//METAWRITE; C; 7; 8; 5
//METAREAD; C; 4
//METAWRITE; A; 1; 2; 3
//METAREAD; A; 4; 5; 6
//METAWRITE; E; 11
//METAREAD; E; 13
//METAWRITE; D; 9
//METAREAD; D; 11
//METAWRITE; F; 13
//METAREAD; F; 1
/////14
